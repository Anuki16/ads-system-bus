
module bus #(
    parameter ADDR_WIDTH = 16,
    parameter DATA_WIDTH = 32
);


endmodule